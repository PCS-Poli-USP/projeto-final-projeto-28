library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity control_unit is
end control_unit;

architecture behaviorial of control_unit is
    
begin

end architecture;