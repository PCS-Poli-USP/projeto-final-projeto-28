library ieee;
use ieee.std_logic_1164.all;

package utils is

    type byte_array is array (integer range <>) of std_logic_vector(7 downto 0);

end utils ;